// my_addition.v  -  ELEC 522 - Fall 2024
// 
// Use these signal names which match the pin constraints .xdc file given
// create a 4 bit unsigned adder using a behavioral description on Zedboard
// add values of sw3, sw2, sw1, sw0 to sw7, sw6, sw5, sw4
// sw0 switch0 is LSB of in_a; sw4 switch4 is LSB of in_b
// display output result in ld4, ld3, ld2, ld1, ld0
// ld4 LED0 is MSB. 


module my_addition (ld4, ld3, ld2, ld1, ld0, sw7, sw6, sw5, sw4, sw3, sw2, sw1, sw0);
	
	// declare port signals
	
	
	
	// declare vectors
	
	
	
	// assign signals to vectors
	
	
	// Add the two four bit numbers; max is 30 or in binary 11110
	
	
  
endmodule
